// RTL (Verilog) generated @ Fri Feb 25 00:20:45 2022 by V3 
//               compiled @ Feb 24 2022 16:36:53
// Internal nets are renamed with prefix "v3_1645719645_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1645719645_0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] v3_1645719645_8;
   reg [2:0] v3_1645719645_9;
   reg [2:0] v3_1645719645_10;
   reg [2:0] v3_1645719645_11;
   reg [1:0] v3_1645719645_12;
   reg [1:0] v3_1645719645_13;
   reg [7:0] v3_1645719645_14;
   reg v3_1645719645_15;
   reg v3_1645719645_16;
   reg [1:0] v3_1645719645_17;
   reg [7:0] v3_1645719645_18;
   reg [2:0] v3_1645719645_19;
   reg [2:0] v3_1645719645_20;
   reg [2:0] v3_1645719645_21;
   reg [2:0] v3_1645719645_22;
   wire [2:0] v3_1645719645_23;
   wire [2:0] v3_1645719645_24;
   wire [2:0] v3_1645719645_25;
   wire [2:0] v3_1645719645_26;
   wire [2:0] v3_1645719645_27;
   wire [2:0] v3_1645719645_28;
   wire [2:0] v3_1645719645_29;
   wire [2:0] v3_1645719645_30;
   wire [2:0] v3_1645719645_31;
   wire [2:0] v3_1645719645_32;
   wire [2:0] v3_1645719645_33;
   wire [2:0] v3_1645719645_34;
   wire [2:0] v3_1645719645_35;
   wire [2:0] v3_1645719645_36;
   wire [2:0] v3_1645719645_37;
   wire v3_1645719645_38;
   wire v3_1645719645_39;
   wire [7:0] v3_1645719645_40;
   wire [7:0] v3_1645719645_41;
   wire v3_1645719645_42;
   wire [1:0] v3_1645719645_43;
   wire [1:0] v3_1645719645_44;
   wire v3_1645719645_45;
   wire [1:0] v3_1645719645_46;
   wire [1:0] v3_1645719645_47;
   wire [2:0] v3_1645719645_48;
   wire [2:0] v3_1645719645_49;
   wire [2:0] v3_1645719645_50;
   wire [2:0] v3_1645719645_51;
   wire [2:0] v3_1645719645_52;
   wire [2:0] v3_1645719645_53;
   wire [2:0] v3_1645719645_54;
   wire v3_1645719645_55;
   wire v3_1645719645_56;
   wire [7:0] v3_1645719645_57;
   wire [7:0] v3_1645719645_58;
   wire v3_1645719645_59;
   wire [1:0] v3_1645719645_60;
   wire [1:0] v3_1645719645_61;
   wire v3_1645719645_62;
   wire [2:0] v3_1645719645_63;
   wire v3_1645719645_64;
   wire [2:0] v3_1645719645_65;
   wire [2:0] v3_1645719645_66;
   wire v3_1645719645_67;
   wire v3_1645719645_68;
   wire v3_1645719645_69;
   wire [2:0] v3_1645719645_70;
   wire v3_1645719645_71;
   wire [2:0] v3_1645719645_72;
   wire [2:0] v3_1645719645_73;
   wire [2:0] v3_1645719645_74;
   wire [2:0] v3_1645719645_75;
   wire [2:0] v3_1645719645_76;
   wire [2:0] v3_1645719645_77;
   wire [2:0] v3_1645719645_78;
   wire [2:0] v3_1645719645_79;
   wire [2:0] v3_1645719645_80;
   wire [2:0] v3_1645719645_81;
   wire [2:0] v3_1645719645_82;
   wire [2:0] v3_1645719645_83;
   wire [2:0] v3_1645719645_84;
   wire [2:0] v3_1645719645_85;
   wire [2:0] v3_1645719645_86;
   wire [2:0] v3_1645719645_87;
   wire [2:0] v3_1645719645_88;
   wire [2:0] v3_1645719645_89;
   wire [2:0] v3_1645719645_90;
   wire v3_1645719645_91;
   wire v3_1645719645_92;
   wire [7:0] v3_1645719645_93;
   wire [7:0] v3_1645719645_94;
   wire [2:0] v3_1645719645_95;
   wire [2:0] v3_1645719645_96;
   wire [2:0] v3_1645719645_97;
   wire [2:0] v3_1645719645_98;
   wire [2:0] v3_1645719645_99;
   wire [2:0] v3_1645719645_100;
   wire [2:0] v3_1645719645_101;
   wire [2:0] v3_1645719645_102;
   wire [2:0] v3_1645719645_103;
   wire [2:0] v3_1645719645_104;
   wire [2:0] v3_1645719645_105;
   wire [2:0] v3_1645719645_106;
   wire [2:0] v3_1645719645_107;
   wire [2:0] v3_1645719645_108;
   wire [2:0] v3_1645719645_109;
   wire [2:0] v3_1645719645_110;
   wire [2:0] v3_1645719645_111;
   wire [2:0] v3_1645719645_112;
   wire [2:0] v3_1645719645_113;
   wire [2:0] v3_1645719645_114;
   wire [2:0] v3_1645719645_115;
   wire [2:0] v3_1645719645_116;
   wire [2:0] v3_1645719645_117;
   wire v3_1645719645_118;
   wire v3_1645719645_119;
   wire [7:0] v3_1645719645_120;
   wire [7:0] v3_1645719645_121;
   wire [2:0] v3_1645719645_122;
   wire [2:0] v3_1645719645_123;
   wire [2:0] v3_1645719645_124;
   wire [2:0] v3_1645719645_125;
   wire [2:0] v3_1645719645_126;
   wire [2:0] v3_1645719645_127;
   wire [2:0] v3_1645719645_128;
   wire [2:0] v3_1645719645_129;
   wire [2:0] v3_1645719645_130;
   wire [2:0] v3_1645719645_131;
   wire [2:0] v3_1645719645_132;
   wire [2:0] v3_1645719645_133;
   wire [2:0] v3_1645719645_134;
   wire [2:0] v3_1645719645_135;
   wire [2:0] v3_1645719645_136;
   wire [2:0] v3_1645719645_137;
   wire [2:0] v3_1645719645_138;
   wire [2:0] v3_1645719645_139;
   wire [2:0] v3_1645719645_140;
   wire [2:0] v3_1645719645_141;
   wire [2:0] v3_1645719645_142;
   wire [2:0] v3_1645719645_143;
   wire [2:0] v3_1645719645_144;
   wire [2:0] v3_1645719645_145;
   wire [2:0] v3_1645719645_146;
   wire [2:0] v3_1645719645_147;
   wire [1:0] v3_1645719645_148;
   wire [1:0] v3_1645719645_149;
   wire [1:0] v3_1645719645_150;
   wire [1:0] v3_1645719645_151;
   wire [1:0] v3_1645719645_152;
   wire [1:0] v3_1645719645_153;
   wire [1:0] v3_1645719645_154;
   wire [1:0] v3_1645719645_155;
   wire [1:0] v3_1645719645_156;
   wire [1:0] v3_1645719645_157;
   wire [1:0] v3_1645719645_158;
   wire [1:0] v3_1645719645_159;
   wire [1:0] v3_1645719645_160;
   wire [1:0] v3_1645719645_161;
   wire [1:0] v3_1645719645_162;
   wire v3_1645719645_163;
   wire v3_1645719645_164;
   wire [1:0] v3_1645719645_165;
   wire [1:0] v3_1645719645_166;
   wire [1:0] v3_1645719645_167;
   wire [1:0] v3_1645719645_168;
   wire [1:0] v3_1645719645_169;
   wire [1:0] v3_1645719645_170;
   wire [1:0] v3_1645719645_171;
   wire [1:0] v3_1645719645_172;
   wire [1:0] v3_1645719645_173;
   wire [1:0] v3_1645719645_174;
   wire [1:0] v3_1645719645_175;
   wire [1:0] v3_1645719645_176;
   wire [1:0] v3_1645719645_177;
   wire [1:0] v3_1645719645_178;
   wire [1:0] v3_1645719645_179;
   wire [1:0] v3_1645719645_180;
   wire [1:0] v3_1645719645_181;
   wire [1:0] v3_1645719645_182;
   wire [1:0] v3_1645719645_183;
   wire [1:0] v3_1645719645_184;
   wire [1:0] v3_1645719645_185;
   wire [1:0] v3_1645719645_186;
   wire [1:0] v3_1645719645_187;
   wire [1:0] v3_1645719645_188;
   wire [7:0] v3_1645719645_189;
   wire [7:0] v3_1645719645_190;
   wire [7:0] v3_1645719645_191;
   wire [7:0] v3_1645719645_192;
   wire [7:0] v3_1645719645_193;
   wire [7:0] v3_1645719645_194;
   wire [7:0] v3_1645719645_195;
   wire [7:0] v3_1645719645_196;
   wire [7:0] v3_1645719645_197;
   wire [7:0] v3_1645719645_198;
   wire [7:0] v3_1645719645_199;
   wire [7:0] v3_1645719645_200;
   wire [7:0] v3_1645719645_201;
   wire [7:0] v3_1645719645_202;
   wire [7:0] v3_1645719645_203;
   wire [7:0] v3_1645719645_204;
   wire [5:0] v3_1645719645_205;
   wire [5:0] v3_1645719645_206;
   wire [7:0] v3_1645719645_207;
   wire [7:0] v3_1645719645_208;
   wire [7:0] v3_1645719645_209;
   wire [7:0] v3_1645719645_210;
   wire [7:0] v3_1645719645_211;
   wire [7:0] v3_1645719645_212;
   wire [7:0] v3_1645719645_213;
   wire [7:0] v3_1645719645_214;
   wire [7:0] v3_1645719645_215;
   wire [7:0] v3_1645719645_216;
   wire [7:0] v3_1645719645_217;
   wire [7:0] v3_1645719645_218;
   wire [7:0] v3_1645719645_219;
   wire [7:0] v3_1645719645_220;
   wire [7:0] v3_1645719645_221;
   wire [7:0] v3_1645719645_222;
   wire [7:0] v3_1645719645_223;
   wire [7:0] v3_1645719645_224;
   wire [7:0] v3_1645719645_225;
   wire [7:0] v3_1645719645_226;
   wire [7:0] v3_1645719645_227;
   wire [7:0] v3_1645719645_228;
   wire [7:0] v3_1645719645_229;
   wire [7:0] v3_1645719645_230;
   wire [7:0] v3_1645719645_231;
   wire [7:0] v3_1645719645_232;
   wire [7:0] v3_1645719645_233;
   wire v3_1645719645_234;
   wire v3_1645719645_235;
   wire v3_1645719645_236;
   wire v3_1645719645_237;
   wire v3_1645719645_238;
   wire v3_1645719645_239;
   wire v3_1645719645_240;
   wire v3_1645719645_241;
   wire v3_1645719645_242;
   wire v3_1645719645_243;
   wire v3_1645719645_244;
   wire v3_1645719645_245;
   wire v3_1645719645_246;
   wire v3_1645719645_247;
   wire v3_1645719645_248;
   wire v3_1645719645_249;
   wire v3_1645719645_250;
   wire v3_1645719645_251;
   wire v3_1645719645_252;
   wire v3_1645719645_253;
   wire v3_1645719645_254;
   wire v3_1645719645_255;
   wire v3_1645719645_256;
   wire [1:0] v3_1645719645_257;
   wire [1:0] v3_1645719645_258;
   wire [1:0] v3_1645719645_259;
   wire [1:0] v3_1645719645_260;
   wire [1:0] v3_1645719645_261;
   wire [1:0] v3_1645719645_262;
   wire [1:0] v3_1645719645_263;
   wire [1:0] v3_1645719645_264;
   wire [1:0] v3_1645719645_265;
   wire [1:0] v3_1645719645_266;
   wire [1:0] v3_1645719645_267;
   wire [1:0] v3_1645719645_268;
   wire [1:0] v3_1645719645_269;
   wire [1:0] v3_1645719645_270;
   wire [1:0] v3_1645719645_271;
   wire [1:0] v3_1645719645_272;
   wire [1:0] v3_1645719645_273;
   wire [1:0] v3_1645719645_274;
   wire [1:0] v3_1645719645_275;
   wire [1:0] v3_1645719645_276;
   wire [1:0] v3_1645719645_277;
   wire [1:0] v3_1645719645_278;
   wire [1:0] v3_1645719645_279;
   wire [1:0] v3_1645719645_280;
   wire [1:0] v3_1645719645_281;
   wire [1:0] v3_1645719645_282;
   wire [1:0] v3_1645719645_283;
   wire [1:0] v3_1645719645_284;
   wire [1:0] v3_1645719645_285;
   wire [1:0] v3_1645719645_286;
   wire [1:0] v3_1645719645_287;
   wire [7:0] v3_1645719645_288;
   wire [7:0] v3_1645719645_289;
   wire [7:0] v3_1645719645_290;
   wire [7:0] v3_1645719645_291;
   wire [7:0] v3_1645719645_292;
   wire [7:0] v3_1645719645_293;
   wire [7:0] v3_1645719645_294;
   wire [7:0] v3_1645719645_295;
   wire [7:0] v3_1645719645_296;
   wire [7:0] v3_1645719645_297;
   wire [7:0] v3_1645719645_298;
   wire [7:0] v3_1645719645_299;
   wire [7:0] v3_1645719645_300;
   wire [7:0] v3_1645719645_301;
   wire [7:0] v3_1645719645_302;
   wire [7:0] v3_1645719645_303;
   wire [7:0] v3_1645719645_304;
   wire [7:0] v3_1645719645_305;
   wire [7:0] v3_1645719645_306;
   wire [7:0] v3_1645719645_307;
   wire [7:0] v3_1645719645_308;
   wire [7:0] v3_1645719645_309;
   wire [7:0] v3_1645719645_310;
   wire [7:0] v3_1645719645_311;
   wire [7:0] v3_1645719645_312;
   wire [7:0] v3_1645719645_313;
   wire [7:0] v3_1645719645_314;
   wire [7:0] v3_1645719645_315;
   wire [7:0] v3_1645719645_316;
   wire [7:0] v3_1645719645_317;
   wire [7:0] v3_1645719645_318;
   wire [7:0] v3_1645719645_319;
   wire [7:0] v3_1645719645_320;
   wire [7:0] v3_1645719645_321;
   wire [7:0] v3_1645719645_322;
   wire [7:0] v3_1645719645_323;
   wire [7:0] v3_1645719645_324;
   wire [7:0] v3_1645719645_325;
   wire [7:0] v3_1645719645_326;
   wire [7:0] v3_1645719645_327;
   wire [7:0] v3_1645719645_328;
   wire [7:0] v3_1645719645_329;
   wire v3_1645719645_330;
   wire [7:0] v3_1645719645_331;
   wire [7:0] v3_1645719645_332;
   wire v3_1645719645_333;
   wire [7:0] v3_1645719645_334;
   wire [7:0] v3_1645719645_335;
   wire v3_1645719645_336;
   wire [7:0] v3_1645719645_337;
   wire [7:0] v3_1645719645_338;
   wire [2:0] v3_1645719645_339;
   wire [2:0] v3_1645719645_340;
   wire [2:0] v3_1645719645_341;
   wire [2:0] v3_1645719645_342;
   wire [2:0] v3_1645719645_343;
   wire [2:0] v3_1645719645_344;
   wire [2:0] v3_1645719645_345;
   wire [2:0] v3_1645719645_346;
   wire [2:0] v3_1645719645_347;
   wire [2:0] v3_1645719645_348;
   wire [2:0] v3_1645719645_349;
   wire [2:0] v3_1645719645_350;
   wire [2:0] v3_1645719645_351;
   wire [2:0] v3_1645719645_352;
   wire [2:0] v3_1645719645_353;
   wire [2:0] v3_1645719645_354;
   wire [2:0] v3_1645719645_355;
   wire [2:0] v3_1645719645_356;
   wire [2:0] v3_1645719645_357;
   wire [2:0] v3_1645719645_358;
   wire [2:0] v3_1645719645_359;
   wire [2:0] v3_1645719645_360;
   wire [2:0] v3_1645719645_361;
   wire [2:0] v3_1645719645_362;
   wire [2:0] v3_1645719645_363;
   wire [2:0] v3_1645719645_364;
   wire [2:0] v3_1645719645_365;
   wire [2:0] v3_1645719645_366;
   wire [2:0] v3_1645719645_367;
   wire [2:0] v3_1645719645_368;
   wire v3_1645719645_369;
   wire [3:0] v3_1645719645_370;
   wire [3:0] v3_1645719645_371;
   wire [3:0] v3_1645719645_372;
   wire [3:0] v3_1645719645_373;
   wire [3:0] v3_1645719645_374;
   wire [3:0] v3_1645719645_375;
   wire [3:0] v3_1645719645_376;
   wire [3:0] v3_1645719645_377;
   wire [3:0] v3_1645719645_378;
   wire [3:0] v3_1645719645_379;
   wire [3:0] v3_1645719645_380;
   wire [2:0] v3_1645719645_381;
   wire [2:0] v3_1645719645_382;
   wire [2:0] v3_1645719645_383;
   wire [2:0] v3_1645719645_384;
   wire [2:0] v3_1645719645_385;
   wire [2:0] v3_1645719645_386;
   wire [2:0] v3_1645719645_387;
   wire [2:0] v3_1645719645_388;
   wire [2:0] v3_1645719645_389;
   wire [2:0] v3_1645719645_390;
   wire [2:0] v3_1645719645_391;
   wire [2:0] v3_1645719645_392;
   wire [2:0] v3_1645719645_393;
   wire [2:0] v3_1645719645_394;
   wire [2:0] v3_1645719645_395;
   wire [2:0] v3_1645719645_396;
   wire [2:0] v3_1645719645_397;
   wire [2:0] v3_1645719645_398;
   wire [2:0] v3_1645719645_399;
   wire [2:0] v3_1645719645_400;
   wire [2:0] v3_1645719645_401;
   wire [2:0] v3_1645719645_402;
   wire [2:0] v3_1645719645_403;
   wire [2:0] v3_1645719645_404;
   wire [2:0] v3_1645719645_405;
   wire [2:0] v3_1645719645_406;
   wire [2:0] v3_1645719645_407;
   wire [2:0] v3_1645719645_408;
   wire [2:0] v3_1645719645_409;
   wire [2:0] v3_1645719645_410;
   wire [2:0] v3_1645719645_411;
   wire [2:0] v3_1645719645_412;
   wire v3_1645719645_413;
   wire [3:0] v3_1645719645_414;
   wire [3:0] v3_1645719645_415;
   wire [3:0] v3_1645719645_416;
   wire [3:0] v3_1645719645_417;
   wire [3:0] v3_1645719645_418;
   wire [3:0] v3_1645719645_419;
   wire [3:0] v3_1645719645_420;
   wire [3:0] v3_1645719645_421;
   wire [3:0] v3_1645719645_422;
   wire [2:0] v3_1645719645_423;
   wire [2:0] v3_1645719645_424;
   wire [2:0] v3_1645719645_425;
   wire [2:0] v3_1645719645_426;
   wire [2:0] v3_1645719645_427;
   wire [2:0] v3_1645719645_428;
   wire [2:0] v3_1645719645_429;
   wire [2:0] v3_1645719645_430;
   wire [2:0] v3_1645719645_431;
   wire [2:0] v3_1645719645_432;
   wire [2:0] v3_1645719645_433;
   wire [2:0] v3_1645719645_434;
   wire [2:0] v3_1645719645_435;
   wire [2:0] v3_1645719645_436;
   wire [2:0] v3_1645719645_437;
   wire [2:0] v3_1645719645_438;
   wire [2:0] v3_1645719645_439;
   wire [2:0] v3_1645719645_440;
   wire [2:0] v3_1645719645_441;
   wire [2:0] v3_1645719645_442;
   wire [2:0] v3_1645719645_443;
   wire [2:0] v3_1645719645_444;
   wire [2:0] v3_1645719645_445;
   wire [2:0] v3_1645719645_446;
   wire [2:0] v3_1645719645_447;
   wire [2:0] v3_1645719645_448;
   wire [2:0] v3_1645719645_449;
   wire [2:0] v3_1645719645_450;
   wire v3_1645719645_451;
   wire [3:0] v3_1645719645_452;
   wire [3:0] v3_1645719645_453;
   wire [3:0] v3_1645719645_454;
   wire [3:0] v3_1645719645_455;
   wire [3:0] v3_1645719645_456;
   wire [3:0] v3_1645719645_457;
   wire [3:0] v3_1645719645_458;
   wire [3:0] v3_1645719645_459;
   wire [3:0] v3_1645719645_460;
   wire [2:0] v3_1645719645_461;
   wire [2:0] v3_1645719645_462;
   wire [2:0] v3_1645719645_463;
   wire [2:0] v3_1645719645_464;
   wire [2:0] v3_1645719645_465;
   wire [2:0] v3_1645719645_466;
   wire [2:0] v3_1645719645_467;
   wire [2:0] v3_1645719645_468;
   wire [2:0] v3_1645719645_469;
   wire [2:0] v3_1645719645_470;
   wire [2:0] v3_1645719645_471;
   wire [2:0] v3_1645719645_472;
   wire [2:0] v3_1645719645_473;
   wire [2:0] v3_1645719645_474;
   wire [2:0] v3_1645719645_475;
   wire [2:0] v3_1645719645_476;
   wire [2:0] v3_1645719645_477;
   wire [2:0] v3_1645719645_478;
   wire [2:0] v3_1645719645_479;
   wire [2:0] v3_1645719645_480;
   wire [2:0] v3_1645719645_481;
   wire [2:0] v3_1645719645_482;
   wire [2:0] v3_1645719645_483;
   wire [2:0] v3_1645719645_484;
   wire [2:0] v3_1645719645_485;
   wire [2:0] v3_1645719645_486;
   wire [2:0] v3_1645719645_487;
   wire [2:0] v3_1645719645_488;
   wire [2:0] v3_1645719645_489;
   wire [2:0] v3_1645719645_490;
   wire v3_1645719645_491;
   wire [3:0] v3_1645719645_492;
   wire [3:0] v3_1645719645_493;
   wire [3:0] v3_1645719645_494;
   wire [3:0] v3_1645719645_495;
   wire [3:0] v3_1645719645_496;
   wire [3:0] v3_1645719645_497;
   wire [3:0] v3_1645719645_498;
   wire [3:0] v3_1645719645_499;
   wire [3:0] v3_1645719645_500;
   wire [2:0] v3_1645719645_501;
   wire [2:0] v3_1645719645_502;
   wire v3_1645719645_503;
   wire v3_1645719645_504;
   wire v3_1645719645_505;
   wire v3_1645719645_506;
   wire v3_1645719645_507;
   wire v3_1645719645_508;
   wire v3_1645719645_509;
   wire v3_1645719645_510;
   wire v3_1645719645_511;
   wire v3_1645719645_512;
   wire v3_1645719645_513;
   wire v3_1645719645_514;
   wire [7:0] v3_1645719645_515;
   wire [7:0] v3_1645719645_516;
   wire [7:0] v3_1645719645_517;
   wire [7:0] v3_1645719645_518;
   wire [7:0] v3_1645719645_519;
   wire [7:0] v3_1645719645_520;
   wire [7:0] v3_1645719645_521;
   wire [7:0] v3_1645719645_522;
   wire [7:0] v3_1645719645_523;
   wire [7:0] v3_1645719645_524;
   wire [4:0] v3_1645719645_525;
   wire [4:0] v3_1645719645_526;
   wire [7:0] v3_1645719645_527;
   wire [7:0] v3_1645719645_528;
   wire [7:0] v3_1645719645_529;
   wire [7:0] v3_1645719645_530;
   wire [7:0] v3_1645719645_531;
   wire [7:0] v3_1645719645_532;
   wire [7:0] v3_1645719645_533;
   wire [7:0] v3_1645719645_534;
   wire [7:0] v3_1645719645_535;
   wire [7:0] v3_1645719645_536;
   wire [7:0] v3_1645719645_537;
   wire [7:0] v3_1645719645_538;
   wire [7:0] v3_1645719645_539;
   wire [7:0] v3_1645719645_540;
   wire [7:0] v3_1645719645_541;
   wire [7:0] v3_1645719645_542;
   wire [7:0] v3_1645719645_543;
   wire [7:0] v3_1645719645_544;
   wire [7:0] v3_1645719645_545;
   wire [7:0] v3_1645719645_546;
   wire [7:0] v3_1645719645_547;
   wire [7:0] v3_1645719645_548;
   wire [7:0] v3_1645719645_549;
   wire v3_1645719645_550;
   wire [2:0] v3_1645719645_551;
   wire [2:0] v3_1645719645_552;
   wire [2:0] v3_1645719645_553;
   wire [2:0] v3_1645719645_554;
   wire [1:0] v3_1645719645_555;
   wire [1:0] v3_1645719645_556;

   // Output Net Declarations
   wire p;
   wire [2:0] coinOutNTD_50;
   wire [2:0] coinOutNTD_10;
   wire [2:0] coinOutNTD_5;
   wire [2:0] coinOutNTD_1;
   wire [1:0] itemTypeOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1645719645_0 = 1'b0; 
   assign v3_1645719645_23 = v3_1645719645_24;
   assign v3_1645719645_24 = v3_1645719645_71 ? v3_1645719645_70 : v3_1645719645_25;
   assign v3_1645719645_25 = v3_1645719645_26;
   assign v3_1645719645_26 = v3_1645719645_69 ? v3_1645719645_65 : v3_1645719645_27;
   assign v3_1645719645_27 = v3_1645719645_64 ? v3_1645719645_63 : v3_1645719645_28;
   assign v3_1645719645_28 = v3_1645719645_62 ? v3_1645719645_33 : v3_1645719645_29;
   assign v3_1645719645_29 = v3_1645719645_59 ? v3_1645719645_48 : v3_1645719645_30;
   assign v3_1645719645_30 = v3_1645719645_45 ? v3_1645719645_33 : v3_1645719645_31;
   assign v3_1645719645_31 = v3_1645719645_42 ? v3_1645719645_33 : v3_1645719645_32;
   assign v3_1645719645_32 = v3_1645719645_39 ? v3_1645719645_34 : v3_1645719645_33;
   assign v3_1645719645_33 = v3_1645719645_8;
   assign v3_1645719645_34 = v3_1645719645_38 ? v3_1645719645_35 : v3_1645719645_33;
   assign v3_1645719645_35 = v3_1645719645_36;
   assign v3_1645719645_36 = v3_1645719645_37;
   assign v3_1645719645_37 = 3'b000; 
   assign v3_1645719645_38 = v3_1645719645_21 == v3_1645719645_36;
   assign v3_1645719645_39 = v3_1645719645_18 >= v3_1645719645_40;
   assign v3_1645719645_40 = v3_1645719645_41;
   assign v3_1645719645_41 = 8'b00000001; 
   assign v3_1645719645_42 = v3_1645719645_17 == v3_1645719645_43;
   assign v3_1645719645_43 = v3_1645719645_44;
   assign v3_1645719645_44 = 2'b10; 
   assign v3_1645719645_45 = v3_1645719645_17 == v3_1645719645_46;
   assign v3_1645719645_46 = v3_1645719645_47;
   assign v3_1645719645_47 = 2'b01; 
   assign v3_1645719645_48 = v3_1645719645_56 ? v3_1645719645_49 : v3_1645719645_33;
   assign v3_1645719645_49 = v3_1645719645_55 ? v3_1645719645_33 : v3_1645719645_50;
   assign v3_1645719645_50 = v3_1645719645_51;
   assign v3_1645719645_51 = v3_1645719645_54;
   assign v3_1645719645_52 = v3_1645719645_53;
   assign v3_1645719645_53 = 3'b001; 
   assign v3_1645719645_54 = v3_1645719645_8 + v3_1645719645_52;
   assign v3_1645719645_55 = v3_1645719645_19 == v3_1645719645_36;
   assign v3_1645719645_56 = v3_1645719645_18 >= v3_1645719645_57;
   assign v3_1645719645_57 = v3_1645719645_58;
   assign v3_1645719645_58 = 8'b00110010; 
   assign v3_1645719645_59 = v3_1645719645_17 == v3_1645719645_60;
   assign v3_1645719645_60 = v3_1645719645_61;
   assign v3_1645719645_61 = 2'b00; 
   assign v3_1645719645_62 = ~v3_1645719645_16;
   assign v3_1645719645_63 = v3_1645719645_36;
   assign v3_1645719645_64 = v3_1645719645_13 == v3_1645719645_60;
   assign v3_1645719645_65 = v3_1645719645_67 ? v3_1645719645_66 : v3_1645719645_33;
   assign v3_1645719645_66 = v3_1645719645_36;
   assign v3_1645719645_67 = ~v3_1645719645_68;
   assign v3_1645719645_68 = itemTypeIn == v3_1645719645_60;
   assign v3_1645719645_69 = v3_1645719645_13 == v3_1645719645_46;
   assign v3_1645719645_70 = v3_1645719645_36;
   assign v3_1645719645_71 = ~reset;
   assign v3_1645719645_72 = 3'b000; 
   assign v3_1645719645_73 = v3_1645719645_74;
   assign v3_1645719645_74 = v3_1645719645_71 ? v3_1645719645_98 : v3_1645719645_75;
   assign v3_1645719645_75 = v3_1645719645_76;
   assign v3_1645719645_76 = v3_1645719645_69 ? v3_1645719645_96 : v3_1645719645_77;
   assign v3_1645719645_77 = v3_1645719645_64 ? v3_1645719645_95 : v3_1645719645_78;
   assign v3_1645719645_78 = v3_1645719645_62 ? v3_1645719645_83 : v3_1645719645_79;
   assign v3_1645719645_79 = v3_1645719645_59 ? v3_1645719645_83 : v3_1645719645_80;
   assign v3_1645719645_80 = v3_1645719645_45 ? v3_1645719645_86 : v3_1645719645_81;
   assign v3_1645719645_81 = v3_1645719645_42 ? v3_1645719645_83 : v3_1645719645_82;
   assign v3_1645719645_82 = v3_1645719645_39 ? v3_1645719645_84 : v3_1645719645_83;
   assign v3_1645719645_83 = v3_1645719645_9;
   assign v3_1645719645_84 = v3_1645719645_38 ? v3_1645719645_85 : v3_1645719645_83;
   assign v3_1645719645_85 = v3_1645719645_36;
   assign v3_1645719645_86 = v3_1645719645_92 ? v3_1645719645_87 : v3_1645719645_83;
   assign v3_1645719645_87 = v3_1645719645_91 ? v3_1645719645_83 : v3_1645719645_88;
   assign v3_1645719645_88 = v3_1645719645_89;
   assign v3_1645719645_89 = v3_1645719645_90;
   assign v3_1645719645_90 = v3_1645719645_9 + v3_1645719645_52;
   assign v3_1645719645_91 = v3_1645719645_20 == v3_1645719645_36;
   assign v3_1645719645_92 = v3_1645719645_18 >= v3_1645719645_93;
   assign v3_1645719645_93 = v3_1645719645_94;
   assign v3_1645719645_94 = 8'b00001010; 
   assign v3_1645719645_95 = v3_1645719645_36;
   assign v3_1645719645_96 = v3_1645719645_67 ? v3_1645719645_97 : v3_1645719645_83;
   assign v3_1645719645_97 = v3_1645719645_36;
   assign v3_1645719645_98 = v3_1645719645_36;
   assign v3_1645719645_99 = 3'b000; 
   assign v3_1645719645_100 = v3_1645719645_101;
   assign v3_1645719645_101 = v3_1645719645_71 ? v3_1645719645_125 : v3_1645719645_102;
   assign v3_1645719645_102 = v3_1645719645_103;
   assign v3_1645719645_103 = v3_1645719645_69 ? v3_1645719645_123 : v3_1645719645_104;
   assign v3_1645719645_104 = v3_1645719645_64 ? v3_1645719645_122 : v3_1645719645_105;
   assign v3_1645719645_105 = v3_1645719645_62 ? v3_1645719645_110 : v3_1645719645_106;
   assign v3_1645719645_106 = v3_1645719645_59 ? v3_1645719645_110 : v3_1645719645_107;
   assign v3_1645719645_107 = v3_1645719645_45 ? v3_1645719645_110 : v3_1645719645_108;
   assign v3_1645719645_108 = v3_1645719645_42 ? v3_1645719645_113 : v3_1645719645_109;
   assign v3_1645719645_109 = v3_1645719645_39 ? v3_1645719645_111 : v3_1645719645_110;
   assign v3_1645719645_110 = v3_1645719645_10;
   assign v3_1645719645_111 = v3_1645719645_38 ? v3_1645719645_112 : v3_1645719645_110;
   assign v3_1645719645_112 = v3_1645719645_36;
   assign v3_1645719645_113 = v3_1645719645_119 ? v3_1645719645_114 : v3_1645719645_110;
   assign v3_1645719645_114 = v3_1645719645_118 ? v3_1645719645_110 : v3_1645719645_115;
   assign v3_1645719645_115 = v3_1645719645_116;
   assign v3_1645719645_116 = v3_1645719645_117;
   assign v3_1645719645_117 = v3_1645719645_10 + v3_1645719645_52;
   assign v3_1645719645_118 = v3_1645719645_22 == v3_1645719645_36;
   assign v3_1645719645_119 = v3_1645719645_18 >= v3_1645719645_120;
   assign v3_1645719645_120 = v3_1645719645_121;
   assign v3_1645719645_121 = 8'b00000101; 
   assign v3_1645719645_122 = v3_1645719645_36;
   assign v3_1645719645_123 = v3_1645719645_67 ? v3_1645719645_124 : v3_1645719645_110;
   assign v3_1645719645_124 = v3_1645719645_36;
   assign v3_1645719645_125 = v3_1645719645_36;
   assign v3_1645719645_126 = 3'b000; 
   assign v3_1645719645_127 = v3_1645719645_128;
   assign v3_1645719645_128 = v3_1645719645_71 ? v3_1645719645_146 : v3_1645719645_129;
   assign v3_1645719645_129 = v3_1645719645_130;
   assign v3_1645719645_130 = v3_1645719645_69 ? v3_1645719645_144 : v3_1645719645_131;
   assign v3_1645719645_131 = v3_1645719645_64 ? v3_1645719645_143 : v3_1645719645_132;
   assign v3_1645719645_132 = v3_1645719645_62 ? v3_1645719645_137 : v3_1645719645_133;
   assign v3_1645719645_133 = v3_1645719645_59 ? v3_1645719645_137 : v3_1645719645_134;
   assign v3_1645719645_134 = v3_1645719645_45 ? v3_1645719645_137 : v3_1645719645_135;
   assign v3_1645719645_135 = v3_1645719645_42 ? v3_1645719645_137 : v3_1645719645_136;
   assign v3_1645719645_136 = v3_1645719645_39 ? v3_1645719645_138 : v3_1645719645_137;
   assign v3_1645719645_137 = v3_1645719645_11;
   assign v3_1645719645_138 = v3_1645719645_38 ? v3_1645719645_142 : v3_1645719645_139;
   assign v3_1645719645_139 = v3_1645719645_140;
   assign v3_1645719645_140 = v3_1645719645_141;
   assign v3_1645719645_141 = v3_1645719645_11 + v3_1645719645_52;
   assign v3_1645719645_142 = v3_1645719645_36;
   assign v3_1645719645_143 = v3_1645719645_36;
   assign v3_1645719645_144 = v3_1645719645_67 ? v3_1645719645_145 : v3_1645719645_137;
   assign v3_1645719645_145 = v3_1645719645_36;
   assign v3_1645719645_146 = v3_1645719645_36;
   assign v3_1645719645_147 = 3'b000; 
   assign v3_1645719645_148 = v3_1645719645_149;
   assign v3_1645719645_149 = v3_1645719645_71 ? v3_1645719645_168 : v3_1645719645_150;
   assign v3_1645719645_150 = v3_1645719645_151;
   assign v3_1645719645_151 = v3_1645719645_69 ? v3_1645719645_166 : v3_1645719645_152;
   assign v3_1645719645_152 = v3_1645719645_64 ? v3_1645719645_165 : v3_1645719645_153;
   assign v3_1645719645_153 = v3_1645719645_62 ? v3_1645719645_161 : v3_1645719645_154;
   assign v3_1645719645_154 = v3_1645719645_59 ? v3_1645719645_158 : v3_1645719645_155;
   assign v3_1645719645_155 = v3_1645719645_45 ? v3_1645719645_158 : v3_1645719645_156;
   assign v3_1645719645_156 = v3_1645719645_42 ? v3_1645719645_158 : v3_1645719645_157;
   assign v3_1645719645_157 = v3_1645719645_39 ? v3_1645719645_159 : v3_1645719645_158;
   assign v3_1645719645_158 = v3_1645719645_12;
   assign v3_1645719645_159 = v3_1645719645_38 ? v3_1645719645_160 : v3_1645719645_158;
   assign v3_1645719645_160 = v3_1645719645_60;
   assign v3_1645719645_161 = v3_1645719645_163 ? v3_1645719645_162 : v3_1645719645_158;
   assign v3_1645719645_162 = v3_1645719645_60;
   assign v3_1645719645_163 = ~v3_1645719645_164;
   assign v3_1645719645_164 = v3_1645719645_14 >= v3_1645719645_18;
   assign v3_1645719645_165 = v3_1645719645_60;
   assign v3_1645719645_166 = v3_1645719645_67 ? v3_1645719645_167 : v3_1645719645_158;
   assign v3_1645719645_167 = itemTypeIn;
   assign v3_1645719645_168 = v3_1645719645_60;
   assign v3_1645719645_169 = 2'b00; 
   assign v3_1645719645_170 = v3_1645719645_171;
   assign v3_1645719645_171 = v3_1645719645_71 ? v3_1645719645_187 : v3_1645719645_172;
   assign v3_1645719645_172 = v3_1645719645_173;
   assign v3_1645719645_173 = v3_1645719645_69 ? v3_1645719645_185 : v3_1645719645_174;
   assign v3_1645719645_174 = v3_1645719645_64 ? v3_1645719645_184 : v3_1645719645_175;
   assign v3_1645719645_175 = v3_1645719645_62 ? v3_1645719645_182 : v3_1645719645_176;
   assign v3_1645719645_176 = v3_1645719645_59 ? v3_1645719645_182 : v3_1645719645_177;
   assign v3_1645719645_177 = v3_1645719645_45 ? v3_1645719645_182 : v3_1645719645_178;
   assign v3_1645719645_178 = v3_1645719645_42 ? v3_1645719645_182 : v3_1645719645_179;
   assign v3_1645719645_179 = v3_1645719645_39 ? v3_1645719645_181 : v3_1645719645_180;
   assign v3_1645719645_180 = v3_1645719645_60;
   assign v3_1645719645_181 = v3_1645719645_38 ? v3_1645719645_183 : v3_1645719645_182;
   assign v3_1645719645_182 = v3_1645719645_13;
   assign v3_1645719645_183 = v3_1645719645_60;
   assign v3_1645719645_184 = v3_1645719645_46;
   assign v3_1645719645_185 = v3_1645719645_67 ? v3_1645719645_186 : v3_1645719645_182;
   assign v3_1645719645_186 = v3_1645719645_43;
   assign v3_1645719645_187 = v3_1645719645_46;
   assign v3_1645719645_188 = 2'b00; 
   assign v3_1645719645_189 = v3_1645719645_190;
   assign v3_1645719645_190 = v3_1645719645_71 ? v3_1645719645_230 : v3_1645719645_191;
   assign v3_1645719645_191 = v3_1645719645_192;
   assign v3_1645719645_192 = v3_1645719645_69 ? v3_1645719645_194 : v3_1645719645_193;
   assign v3_1645719645_193 = v3_1645719645_14;
   assign v3_1645719645_194 = v3_1645719645_67 ? v3_1645719645_195 : v3_1645719645_193;
   assign v3_1645719645_195 = v3_1645719645_196;
   assign v3_1645719645_196 = v3_1645719645_229;
   assign v3_1645719645_197 = v3_1645719645_198;
   assign v3_1645719645_198 = v3_1645719645_222;
   assign v3_1645719645_199 = v3_1645719645_200;
   assign v3_1645719645_200 = v3_1645719645_215;
   assign v3_1645719645_201 = v3_1645719645_202;
   assign v3_1645719645_202 = v3_1645719645_208;
   assign v3_1645719645_203 = v3_1645719645_204;
   assign v3_1645719645_204 = v3_1645719645_207;
   assign v3_1645719645_205 = v3_1645719645_206;
   assign v3_1645719645_206 = 6'b000000; 
   assign v3_1645719645_207 = {v3_1645719645_205, coinInNTD_50};
   assign v3_1645719645_208 = v3_1645719645_57 * v3_1645719645_203;
   assign v3_1645719645_209 = v3_1645719645_210;
   assign v3_1645719645_210 = v3_1645719645_214;
   assign v3_1645719645_211 = v3_1645719645_212;
   assign v3_1645719645_212 = v3_1645719645_213;
   assign v3_1645719645_213 = {v3_1645719645_205, coinInNTD_10};
   assign v3_1645719645_214 = v3_1645719645_93 * v3_1645719645_211;
   assign v3_1645719645_215 = v3_1645719645_201 + v3_1645719645_209;
   assign v3_1645719645_216 = v3_1645719645_217;
   assign v3_1645719645_217 = v3_1645719645_221;
   assign v3_1645719645_218 = v3_1645719645_219;
   assign v3_1645719645_219 = v3_1645719645_220;
   assign v3_1645719645_220 = {v3_1645719645_205, coinInNTD_5};
   assign v3_1645719645_221 = v3_1645719645_120 * v3_1645719645_218;
   assign v3_1645719645_222 = v3_1645719645_199 + v3_1645719645_216;
   assign v3_1645719645_223 = v3_1645719645_224;
   assign v3_1645719645_224 = v3_1645719645_228;
   assign v3_1645719645_225 = v3_1645719645_226;
   assign v3_1645719645_226 = v3_1645719645_227;
   assign v3_1645719645_227 = {v3_1645719645_205, coinInNTD_1};
   assign v3_1645719645_228 = v3_1645719645_40 * v3_1645719645_225;
   assign v3_1645719645_229 = v3_1645719645_197 + v3_1645719645_223;
   assign v3_1645719645_230 = v3_1645719645_231;
   assign v3_1645719645_231 = v3_1645719645_232;
   assign v3_1645719645_232 = 8'b00000000; 
   assign v3_1645719645_233 = 8'b00000000; 
   assign v3_1645719645_234 = v3_1645719645_235;
   assign v3_1645719645_235 = v3_1645719645_71 ? v3_1645719645_237 : v3_1645719645_236;
   assign v3_1645719645_236 = v3_1645719645_15;
   assign v3_1645719645_237 = v3_1645719645_238;
   assign v3_1645719645_238 = v3_1645719645_239;
   assign v3_1645719645_239 = 1'b1; 
   assign v3_1645719645_240 = 1'b0; 
   assign v3_1645719645_241 = v3_1645719645_242;
   assign v3_1645719645_242 = v3_1645719645_71 ? v3_1645719645_255 : v3_1645719645_243;
   assign v3_1645719645_243 = v3_1645719645_244;
   assign v3_1645719645_244 = v3_1645719645_69 ? v3_1645719645_251 : v3_1645719645_245;
   assign v3_1645719645_245 = v3_1645719645_64 ? v3_1645719645_247 : v3_1645719645_246;
   assign v3_1645719645_246 = v3_1645719645_62 ? v3_1645719645_248 : v3_1645719645_247;
   assign v3_1645719645_247 = v3_1645719645_16;
   assign v3_1645719645_248 = v3_1645719645_163 ? v3_1645719645_250 : v3_1645719645_249;
   assign v3_1645719645_249 = v3_1645719645_238;
   assign v3_1645719645_250 = v3_1645719645_238;
   assign v3_1645719645_251 = v3_1645719645_67 ? v3_1645719645_252 : v3_1645719645_247;
   assign v3_1645719645_252 = v3_1645719645_253;
   assign v3_1645719645_253 = v3_1645719645_254;
   assign v3_1645719645_254 = 1'b0; 
   assign v3_1645719645_255 = v3_1645719645_253;
   assign v3_1645719645_256 = 1'b0; 
   assign v3_1645719645_257 = v3_1645719645_258;
   assign v3_1645719645_258 = v3_1645719645_71 ? v3_1645719645_286 : v3_1645719645_259;
   assign v3_1645719645_259 = v3_1645719645_260;
   assign v3_1645719645_260 = v3_1645719645_69 ? v3_1645719645_284 : v3_1645719645_261;
   assign v3_1645719645_261 = v3_1645719645_64 ? v3_1645719645_267 : v3_1645719645_262;
   assign v3_1645719645_262 = v3_1645719645_62 ? v3_1645719645_267 : v3_1645719645_263;
   assign v3_1645719645_263 = v3_1645719645_59 ? v3_1645719645_280 : v3_1645719645_264;
   assign v3_1645719645_264 = v3_1645719645_45 ? v3_1645719645_276 : v3_1645719645_265;
   assign v3_1645719645_265 = v3_1645719645_42 ? v3_1645719645_270 : v3_1645719645_266;
   assign v3_1645719645_266 = v3_1645719645_39 ? v3_1645719645_268 : v3_1645719645_267;
   assign v3_1645719645_267 = v3_1645719645_17;
   assign v3_1645719645_268 = v3_1645719645_38 ? v3_1645719645_269 : v3_1645719645_267;
   assign v3_1645719645_269 = v3_1645719645_60;
   assign v3_1645719645_270 = v3_1645719645_119 ? v3_1645719645_274 : v3_1645719645_271;
   assign v3_1645719645_271 = v3_1645719645_272;
   assign v3_1645719645_272 = v3_1645719645_273;
   assign v3_1645719645_273 = 2'b11; 
   assign v3_1645719645_274 = v3_1645719645_118 ? v3_1645719645_275 : v3_1645719645_267;
   assign v3_1645719645_275 = v3_1645719645_272;
   assign v3_1645719645_276 = v3_1645719645_92 ? v3_1645719645_278 : v3_1645719645_277;
   assign v3_1645719645_277 = v3_1645719645_43;
   assign v3_1645719645_278 = v3_1645719645_91 ? v3_1645719645_279 : v3_1645719645_267;
   assign v3_1645719645_279 = v3_1645719645_43;
   assign v3_1645719645_280 = v3_1645719645_56 ? v3_1645719645_282 : v3_1645719645_281;
   assign v3_1645719645_281 = v3_1645719645_46;
   assign v3_1645719645_282 = v3_1645719645_55 ? v3_1645719645_283 : v3_1645719645_267;
   assign v3_1645719645_283 = v3_1645719645_46;
   assign v3_1645719645_284 = v3_1645719645_67 ? v3_1645719645_285 : v3_1645719645_267;
   assign v3_1645719645_285 = v3_1645719645_60;
   assign v3_1645719645_286 = v3_1645719645_60;
   assign v3_1645719645_287 = 2'b00; 
   assign v3_1645719645_288 = v3_1645719645_289;
   assign v3_1645719645_289 = v3_1645719645_71 ? v3_1645719645_337 : v3_1645719645_290;
   assign v3_1645719645_290 = v3_1645719645_291;
   assign v3_1645719645_291 = v3_1645719645_69 ? v3_1645719645_324 : v3_1645719645_292;
   assign v3_1645719645_292 = v3_1645719645_64 ? v3_1645719645_298 : v3_1645719645_293;
   assign v3_1645719645_293 = v3_1645719645_62 ? v3_1645719645_319 : v3_1645719645_294;
   assign v3_1645719645_294 = v3_1645719645_59 ? v3_1645719645_314 : v3_1645719645_295;
   assign v3_1645719645_295 = v3_1645719645_45 ? v3_1645719645_309 : v3_1645719645_296;
   assign v3_1645719645_296 = v3_1645719645_42 ? v3_1645719645_304 : v3_1645719645_297;
   assign v3_1645719645_297 = v3_1645719645_39 ? v3_1645719645_299 : v3_1645719645_298;
   assign v3_1645719645_298 = v3_1645719645_18;
   assign v3_1645719645_299 = v3_1645719645_38 ? v3_1645719645_303 : v3_1645719645_300;
   assign v3_1645719645_300 = v3_1645719645_301;
   assign v3_1645719645_301 = v3_1645719645_302;
   assign v3_1645719645_302 = v3_1645719645_18 - v3_1645719645_40;
   assign v3_1645719645_303 = v3_1645719645_14;
   assign v3_1645719645_304 = v3_1645719645_119 ? v3_1645719645_305 : v3_1645719645_298;
   assign v3_1645719645_305 = v3_1645719645_118 ? v3_1645719645_298 : v3_1645719645_306;
   assign v3_1645719645_306 = v3_1645719645_307;
   assign v3_1645719645_307 = v3_1645719645_308;
   assign v3_1645719645_308 = v3_1645719645_18 - v3_1645719645_120;
   assign v3_1645719645_309 = v3_1645719645_92 ? v3_1645719645_310 : v3_1645719645_298;
   assign v3_1645719645_310 = v3_1645719645_91 ? v3_1645719645_298 : v3_1645719645_311;
   assign v3_1645719645_311 = v3_1645719645_312;
   assign v3_1645719645_312 = v3_1645719645_313;
   assign v3_1645719645_313 = v3_1645719645_18 - v3_1645719645_93;
   assign v3_1645719645_314 = v3_1645719645_56 ? v3_1645719645_315 : v3_1645719645_298;
   assign v3_1645719645_315 = v3_1645719645_55 ? v3_1645719645_298 : v3_1645719645_316;
   assign v3_1645719645_316 = v3_1645719645_317;
   assign v3_1645719645_317 = v3_1645719645_318;
   assign v3_1645719645_318 = v3_1645719645_18 - v3_1645719645_57;
   assign v3_1645719645_319 = v3_1645719645_163 ? v3_1645719645_323 : v3_1645719645_320;
   assign v3_1645719645_320 = v3_1645719645_321;
   assign v3_1645719645_321 = v3_1645719645_322;
   assign v3_1645719645_322 = v3_1645719645_14 - v3_1645719645_18;
   assign v3_1645719645_323 = v3_1645719645_14;
   assign v3_1645719645_324 = v3_1645719645_67 ? v3_1645719645_325 : v3_1645719645_298;
   assign v3_1645719645_325 = v3_1645719645_336 ? v3_1645719645_334 : v3_1645719645_326;
   assign v3_1645719645_326 = v3_1645719645_333 ? v3_1645719645_331 : v3_1645719645_327;
   assign v3_1645719645_327 = v3_1645719645_330 ? v3_1645719645_328 : v3_1645719645_231;
   assign v3_1645719645_328 = v3_1645719645_329;
   assign v3_1645719645_329 = 8'b00010110; 
   assign v3_1645719645_330 = itemTypeIn == v3_1645719645_272;
   assign v3_1645719645_331 = v3_1645719645_332;
   assign v3_1645719645_332 = 8'b00001111; 
   assign v3_1645719645_333 = itemTypeIn == v3_1645719645_43;
   assign v3_1645719645_334 = v3_1645719645_335;
   assign v3_1645719645_335 = 8'b00001000; 
   assign v3_1645719645_336 = itemTypeIn == v3_1645719645_46;
   assign v3_1645719645_337 = v3_1645719645_231;
   assign v3_1645719645_338 = 8'b00000000; 
   assign v3_1645719645_339 = v3_1645719645_340;
   assign v3_1645719645_340 = v3_1645719645_71 ? v3_1645719645_381 : v3_1645719645_341;
   assign v3_1645719645_341 = v3_1645719645_342;
   assign v3_1645719645_342 = v3_1645719645_69 ? v3_1645719645_359 : v3_1645719645_343;
   assign v3_1645719645_343 = v3_1645719645_64 ? v3_1645719645_349 : v3_1645719645_344;
   assign v3_1645719645_344 = v3_1645719645_62 ? v3_1645719645_349 : v3_1645719645_345;
   assign v3_1645719645_345 = v3_1645719645_59 ? v3_1645719645_354 : v3_1645719645_346;
   assign v3_1645719645_346 = v3_1645719645_45 ? v3_1645719645_349 : v3_1645719645_347;
   assign v3_1645719645_347 = v3_1645719645_42 ? v3_1645719645_349 : v3_1645719645_348;
   assign v3_1645719645_348 = v3_1645719645_39 ? v3_1645719645_350 : v3_1645719645_349;
   assign v3_1645719645_349 = v3_1645719645_19;
   assign v3_1645719645_350 = v3_1645719645_38 ? v3_1645719645_351 : v3_1645719645_349;
   assign v3_1645719645_351 = v3_1645719645_352;
   assign v3_1645719645_352 = v3_1645719645_353;
   assign v3_1645719645_353 = v3_1645719645_19 + v3_1645719645_8;
   assign v3_1645719645_354 = v3_1645719645_56 ? v3_1645719645_355 : v3_1645719645_349;
   assign v3_1645719645_355 = v3_1645719645_55 ? v3_1645719645_349 : v3_1645719645_356;
   assign v3_1645719645_356 = v3_1645719645_357;
   assign v3_1645719645_357 = v3_1645719645_358;
   assign v3_1645719645_358 = v3_1645719645_19 - v3_1645719645_52;
   assign v3_1645719645_359 = v3_1645719645_67 ? v3_1645719645_360 : v3_1645719645_349;
   assign v3_1645719645_360 = v3_1645719645_369 ? v3_1645719645_367 : v3_1645719645_361;
   assign v3_1645719645_361 = v3_1645719645_362;
   assign v3_1645719645_362 = v3_1645719645_366;
   assign v3_1645719645_363 = v3_1645719645_364;
   assign v3_1645719645_364 = v3_1645719645_365;
   assign v3_1645719645_365 = {v3_1645719645_253, coinInNTD_50};
   assign v3_1645719645_366 = v3_1645719645_19 + v3_1645719645_363;
   assign v3_1645719645_367 = v3_1645719645_368;
   assign v3_1645719645_368 = 3'b111; 
   assign v3_1645719645_369 = v3_1645719645_370 >= v3_1645719645_379;
   assign v3_1645719645_370 = v3_1645719645_371;
   assign v3_1645719645_371 = v3_1645719645_378;
   assign v3_1645719645_372 = v3_1645719645_373;
   assign v3_1645719645_373 = v3_1645719645_374;
   assign v3_1645719645_374 = {v3_1645719645_253, v3_1645719645_19};
   assign v3_1645719645_375 = v3_1645719645_376;
   assign v3_1645719645_376 = v3_1645719645_377;
   assign v3_1645719645_377 = {v3_1645719645_60, coinInNTD_50};
   assign v3_1645719645_378 = v3_1645719645_372 + v3_1645719645_375;
   assign v3_1645719645_379 = v3_1645719645_380;
   assign v3_1645719645_380 = 4'b0111; 
   assign v3_1645719645_381 = v3_1645719645_382;
   assign v3_1645719645_382 = v3_1645719645_383;
   assign v3_1645719645_383 = 3'b010; 
   assign v3_1645719645_384 = 3'b000; 
   assign v3_1645719645_385 = v3_1645719645_386;
   assign v3_1645719645_386 = v3_1645719645_71 ? v3_1645719645_423 : v3_1645719645_387;
   assign v3_1645719645_387 = v3_1645719645_388;
   assign v3_1645719645_388 = v3_1645719645_69 ? v3_1645719645_405 : v3_1645719645_389;
   assign v3_1645719645_389 = v3_1645719645_64 ? v3_1645719645_395 : v3_1645719645_390;
   assign v3_1645719645_390 = v3_1645719645_62 ? v3_1645719645_395 : v3_1645719645_391;
   assign v3_1645719645_391 = v3_1645719645_59 ? v3_1645719645_395 : v3_1645719645_392;
   assign v3_1645719645_392 = v3_1645719645_45 ? v3_1645719645_400 : v3_1645719645_393;
   assign v3_1645719645_393 = v3_1645719645_42 ? v3_1645719645_395 : v3_1645719645_394;
   assign v3_1645719645_394 = v3_1645719645_39 ? v3_1645719645_396 : v3_1645719645_395;
   assign v3_1645719645_395 = v3_1645719645_20;
   assign v3_1645719645_396 = v3_1645719645_38 ? v3_1645719645_397 : v3_1645719645_395;
   assign v3_1645719645_397 = v3_1645719645_398;
   assign v3_1645719645_398 = v3_1645719645_399;
   assign v3_1645719645_399 = v3_1645719645_20 + v3_1645719645_9;
   assign v3_1645719645_400 = v3_1645719645_92 ? v3_1645719645_401 : v3_1645719645_395;
   assign v3_1645719645_401 = v3_1645719645_91 ? v3_1645719645_395 : v3_1645719645_402;
   assign v3_1645719645_402 = v3_1645719645_403;
   assign v3_1645719645_403 = v3_1645719645_404;
   assign v3_1645719645_404 = v3_1645719645_20 - v3_1645719645_52;
   assign v3_1645719645_405 = v3_1645719645_67 ? v3_1645719645_406 : v3_1645719645_395;
   assign v3_1645719645_406 = v3_1645719645_413 ? v3_1645719645_367 : v3_1645719645_407;
   assign v3_1645719645_407 = v3_1645719645_408;
   assign v3_1645719645_408 = v3_1645719645_412;
   assign v3_1645719645_409 = v3_1645719645_410;
   assign v3_1645719645_410 = v3_1645719645_411;
   assign v3_1645719645_411 = {v3_1645719645_253, coinInNTD_10};
   assign v3_1645719645_412 = v3_1645719645_20 + v3_1645719645_409;
   assign v3_1645719645_413 = v3_1645719645_414 >= v3_1645719645_379;
   assign v3_1645719645_414 = v3_1645719645_415;
   assign v3_1645719645_415 = v3_1645719645_422;
   assign v3_1645719645_416 = v3_1645719645_417;
   assign v3_1645719645_417 = v3_1645719645_418;
   assign v3_1645719645_418 = {v3_1645719645_253, v3_1645719645_20};
   assign v3_1645719645_419 = v3_1645719645_420;
   assign v3_1645719645_420 = v3_1645719645_421;
   assign v3_1645719645_421 = {v3_1645719645_60, coinInNTD_10};
   assign v3_1645719645_422 = v3_1645719645_416 + v3_1645719645_419;
   assign v3_1645719645_423 = v3_1645719645_382;
   assign v3_1645719645_424 = 3'b000; 
   assign v3_1645719645_425 = v3_1645719645_426;
   assign v3_1645719645_426 = v3_1645719645_71 ? v3_1645719645_461 : v3_1645719645_427;
   assign v3_1645719645_427 = v3_1645719645_428;
   assign v3_1645719645_428 = v3_1645719645_69 ? v3_1645719645_443 : v3_1645719645_429;
   assign v3_1645719645_429 = v3_1645719645_64 ? v3_1645719645_435 : v3_1645719645_430;
   assign v3_1645719645_430 = v3_1645719645_62 ? v3_1645719645_435 : v3_1645719645_431;
   assign v3_1645719645_431 = v3_1645719645_59 ? v3_1645719645_435 : v3_1645719645_432;
   assign v3_1645719645_432 = v3_1645719645_45 ? v3_1645719645_435 : v3_1645719645_433;
   assign v3_1645719645_433 = v3_1645719645_42 ? v3_1645719645_435 : v3_1645719645_434;
   assign v3_1645719645_434 = v3_1645719645_39 ? v3_1645719645_436 : v3_1645719645_435;
   assign v3_1645719645_435 = v3_1645719645_21;
   assign v3_1645719645_436 = v3_1645719645_38 ? v3_1645719645_440 : v3_1645719645_437;
   assign v3_1645719645_437 = v3_1645719645_438;
   assign v3_1645719645_438 = v3_1645719645_439;
   assign v3_1645719645_439 = v3_1645719645_21 - v3_1645719645_52;
   assign v3_1645719645_440 = v3_1645719645_441;
   assign v3_1645719645_441 = v3_1645719645_442;
   assign v3_1645719645_442 = v3_1645719645_21 + v3_1645719645_11;
   assign v3_1645719645_443 = v3_1645719645_67 ? v3_1645719645_444 : v3_1645719645_435;
   assign v3_1645719645_444 = v3_1645719645_451 ? v3_1645719645_367 : v3_1645719645_445;
   assign v3_1645719645_445 = v3_1645719645_446;
   assign v3_1645719645_446 = v3_1645719645_450;
   assign v3_1645719645_447 = v3_1645719645_448;
   assign v3_1645719645_448 = v3_1645719645_449;
   assign v3_1645719645_449 = {v3_1645719645_253, coinInNTD_1};
   assign v3_1645719645_450 = v3_1645719645_21 + v3_1645719645_447;
   assign v3_1645719645_451 = v3_1645719645_452 >= v3_1645719645_379;
   assign v3_1645719645_452 = v3_1645719645_453;
   assign v3_1645719645_453 = v3_1645719645_460;
   assign v3_1645719645_454 = v3_1645719645_455;
   assign v3_1645719645_455 = v3_1645719645_456;
   assign v3_1645719645_456 = {v3_1645719645_253, v3_1645719645_21};
   assign v3_1645719645_457 = v3_1645719645_458;
   assign v3_1645719645_458 = v3_1645719645_459;
   assign v3_1645719645_459 = {v3_1645719645_60, coinInNTD_1};
   assign v3_1645719645_460 = v3_1645719645_454 + v3_1645719645_457;
   assign v3_1645719645_461 = v3_1645719645_382;
   assign v3_1645719645_462 = 3'b000; 
   assign v3_1645719645_463 = v3_1645719645_464;
   assign v3_1645719645_464 = v3_1645719645_71 ? v3_1645719645_501 : v3_1645719645_465;
   assign v3_1645719645_465 = v3_1645719645_466;
   assign v3_1645719645_466 = v3_1645719645_69 ? v3_1645719645_483 : v3_1645719645_467;
   assign v3_1645719645_467 = v3_1645719645_64 ? v3_1645719645_473 : v3_1645719645_468;
   assign v3_1645719645_468 = v3_1645719645_62 ? v3_1645719645_473 : v3_1645719645_469;
   assign v3_1645719645_469 = v3_1645719645_59 ? v3_1645719645_473 : v3_1645719645_470;
   assign v3_1645719645_470 = v3_1645719645_45 ? v3_1645719645_473 : v3_1645719645_471;
   assign v3_1645719645_471 = v3_1645719645_42 ? v3_1645719645_478 : v3_1645719645_472;
   assign v3_1645719645_472 = v3_1645719645_39 ? v3_1645719645_474 : v3_1645719645_473;
   assign v3_1645719645_473 = v3_1645719645_22;
   assign v3_1645719645_474 = v3_1645719645_38 ? v3_1645719645_475 : v3_1645719645_473;
   assign v3_1645719645_475 = v3_1645719645_476;
   assign v3_1645719645_476 = v3_1645719645_477;
   assign v3_1645719645_477 = v3_1645719645_22 + v3_1645719645_10;
   assign v3_1645719645_478 = v3_1645719645_119 ? v3_1645719645_479 : v3_1645719645_473;
   assign v3_1645719645_479 = v3_1645719645_118 ? v3_1645719645_473 : v3_1645719645_480;
   assign v3_1645719645_480 = v3_1645719645_481;
   assign v3_1645719645_481 = v3_1645719645_482;
   assign v3_1645719645_482 = v3_1645719645_22 - v3_1645719645_52;
   assign v3_1645719645_483 = v3_1645719645_67 ? v3_1645719645_484 : v3_1645719645_473;
   assign v3_1645719645_484 = v3_1645719645_491 ? v3_1645719645_367 : v3_1645719645_485;
   assign v3_1645719645_485 = v3_1645719645_486;
   assign v3_1645719645_486 = v3_1645719645_490;
   assign v3_1645719645_487 = v3_1645719645_488;
   assign v3_1645719645_488 = v3_1645719645_489;
   assign v3_1645719645_489 = {v3_1645719645_253, coinInNTD_5};
   assign v3_1645719645_490 = v3_1645719645_22 + v3_1645719645_487;
   assign v3_1645719645_491 = v3_1645719645_492 >= v3_1645719645_379;
   assign v3_1645719645_492 = v3_1645719645_493;
   assign v3_1645719645_493 = v3_1645719645_500;
   assign v3_1645719645_494 = v3_1645719645_495;
   assign v3_1645719645_495 = v3_1645719645_496;
   assign v3_1645719645_496 = {v3_1645719645_253, v3_1645719645_22};
   assign v3_1645719645_497 = v3_1645719645_498;
   assign v3_1645719645_498 = v3_1645719645_499;
   assign v3_1645719645_499 = {v3_1645719645_60, coinInNTD_5};
   assign v3_1645719645_500 = v3_1645719645_494 + v3_1645719645_497;
   assign v3_1645719645_501 = v3_1645719645_382;
   assign v3_1645719645_502 = 3'b000; 
   assign v3_1645719645_503 = v3_1645719645_504;
   assign v3_1645719645_504 = v3_1645719645_505;
   assign v3_1645719645_505 = v3_1645719645_550;
   assign v3_1645719645_506 = v3_1645719645_507;
   assign v3_1645719645_507 = v3_1645719645_512;
   assign v3_1645719645_508 = v3_1645719645_509;
   assign v3_1645719645_509 = v3_1645719645_510;
   assign v3_1645719645_510 = v3_1645719645_15 & v3_1645719645_64;
   assign v3_1645719645_511 = v3_1645719645_12 == v3_1645719645_60;
   assign v3_1645719645_512 = v3_1645719645_508 & v3_1645719645_511;
   assign v3_1645719645_513 = ~v3_1645719645_514;
   assign v3_1645719645_514 = v3_1645719645_515 == v3_1645719645_14;
   assign v3_1645719645_515 = v3_1645719645_516;
   assign v3_1645719645_516 = v3_1645719645_549;
   assign v3_1645719645_517 = v3_1645719645_518;
   assign v3_1645719645_518 = v3_1645719645_542;
   assign v3_1645719645_519 = v3_1645719645_520;
   assign v3_1645719645_520 = v3_1645719645_535;
   assign v3_1645719645_521 = v3_1645719645_522;
   assign v3_1645719645_522 = v3_1645719645_528;
   assign v3_1645719645_523 = v3_1645719645_524;
   assign v3_1645719645_524 = v3_1645719645_527;
   assign v3_1645719645_525 = v3_1645719645_526;
   assign v3_1645719645_526 = 5'b00000; 
   assign v3_1645719645_527 = {v3_1645719645_525, v3_1645719645_8};
   assign v3_1645719645_528 = v3_1645719645_57 * v3_1645719645_523;
   assign v3_1645719645_529 = v3_1645719645_530;
   assign v3_1645719645_530 = v3_1645719645_534;
   assign v3_1645719645_531 = v3_1645719645_532;
   assign v3_1645719645_532 = v3_1645719645_533;
   assign v3_1645719645_533 = {v3_1645719645_525, v3_1645719645_9};
   assign v3_1645719645_534 = v3_1645719645_93 * v3_1645719645_531;
   assign v3_1645719645_535 = v3_1645719645_521 + v3_1645719645_529;
   assign v3_1645719645_536 = v3_1645719645_537;
   assign v3_1645719645_537 = v3_1645719645_541;
   assign v3_1645719645_538 = v3_1645719645_539;
   assign v3_1645719645_539 = v3_1645719645_540;
   assign v3_1645719645_540 = {v3_1645719645_525, v3_1645719645_10};
   assign v3_1645719645_541 = v3_1645719645_120 * v3_1645719645_538;
   assign v3_1645719645_542 = v3_1645719645_519 + v3_1645719645_536;
   assign v3_1645719645_543 = v3_1645719645_544;
   assign v3_1645719645_544 = v3_1645719645_548;
   assign v3_1645719645_545 = v3_1645719645_546;
   assign v3_1645719645_546 = v3_1645719645_547;
   assign v3_1645719645_547 = {v3_1645719645_525, v3_1645719645_11};
   assign v3_1645719645_548 = v3_1645719645_40 * v3_1645719645_545;
   assign v3_1645719645_549 = v3_1645719645_517 + v3_1645719645_543;
   assign v3_1645719645_550 = v3_1645719645_506 & v3_1645719645_513;
   assign v3_1645719645_551 = v3_1645719645_8;
   assign v3_1645719645_552 = v3_1645719645_9;
   assign v3_1645719645_553 = v3_1645719645_10;
   assign v3_1645719645_554 = v3_1645719645_11;
   assign v3_1645719645_555 = v3_1645719645_12;
   assign v3_1645719645_556 = v3_1645719645_13;

   // Output Net Assignments
   assign p = v3_1645719645_503;
   assign coinOutNTD_50 = v3_1645719645_551;
   assign coinOutNTD_10 = v3_1645719645_552;
   assign coinOutNTD_5 = v3_1645719645_553;
   assign coinOutNTD_1 = v3_1645719645_554;
   assign itemTypeOut = v3_1645719645_555;
   assign serviceTypeOut = v3_1645719645_556;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1645719645_8 <= v3_1645719645_23;
      v3_1645719645_9 <= v3_1645719645_73;
      v3_1645719645_10 <= v3_1645719645_100;
      v3_1645719645_11 <= v3_1645719645_127;
      v3_1645719645_12 <= v3_1645719645_148;
      v3_1645719645_13 <= v3_1645719645_170;
      v3_1645719645_14 <= v3_1645719645_189;
      v3_1645719645_15 <= v3_1645719645_234;
      v3_1645719645_16 <= v3_1645719645_241;
      v3_1645719645_17 <= v3_1645719645_257;
      v3_1645719645_18 <= v3_1645719645_288;
      v3_1645719645_19 <= v3_1645719645_339;
      v3_1645719645_20 <= v3_1645719645_385;
      v3_1645719645_21 <= v3_1645719645_425;
      v3_1645719645_22 <= v3_1645719645_463;
   end
endmodule
